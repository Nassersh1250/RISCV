`timescale 1ns / 1ps

module Data_memory(
    input logic clk,resetn,memwrite,
    input logic [31:0]addr, wdata,
    output logic [31:0] rdata
    );
    
    always@(*) begin
        rdata
endmodule
